`ifndef rhlib__sv
`define rhlib__sv

package Rhlib;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "rhTypes.svh"
	`include "rhResetTransBase.svh"
	`include "rhMonitorBase.svh"
	`include "rhDriverBase.svh"
endpackage

`endif
