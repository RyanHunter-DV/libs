`ifndef RHGpVipPkg__sv
`define RHGpVipPkg__sv

`include "uvm_macros.svh"
`include "GpvInterface.sv"
package RHGpVipPkg;

	import uvm_pkg::*;

	`include "GpvTypes.svh"
	`include "GpvSeqItem.svh"
	`include "GpvDriveVectors.svh"
	`include "GpvInterfaceMap.svh"
	`include "GpvDriveObject.svh"
	`include "GpvProtocoolBase.svh"
	`include "GpvDriver.svh"
	`include "GpvSeqr.svh"
	`include "GpvAgent.svh"

endpackage

`endif
