`ifndef VipBaseTypes__svh
`define VipBaseTypes__svh


typedef enum {
	resetActive,
	resetInActive,
	resetUnknown
}VipResetStatus;

`endif
