typedef enum bit {
	false = 1'b0,
	true  = 1'b1
}bool;
