`ifndef rh_stdint__svh
`define rh_stdint__svh

typedef int unsigned uint32_t;



`endif
