`ifndef RHVipBase__sv
`define RHVipBase__sv

package RHVipBase; // {

	`include "uvm_macros.svh"
	import uvm_pkg::*;


	`include "VipBaseTypes.svh"
	`include "VipResetTrans.svh"
	`include "VipEnvBase.svh"
	`include "VipMonitorBase.svh"
	`include "VipDriverBase.svh"
	`include "VipResetHandler.svh"
	`include "VipAgentBase.svh"



endpackage // }

`endif
