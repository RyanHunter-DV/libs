`ifndef rhGpv__sv
`define rhGpv__sv

`include "rhGpvIf.sv"
package RhGpv;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "rhlib.sv"
	import RhLib::*;
	`include "rhGpvTypes.svh"
	
	`include "rhGpvInterfaceControl.svh"
	`include "rhGpvConfig.svh"
	`include "rhGpvDriveObject.svh"
	`include "rhGpvProtocolBase.svh"
	
	`include "rhGpvDriver.svh"
	`include "rhGpvMonitor.svh"
	`include "rhGpvAgent.svh"
endpackage

`endif
