`ifndef GpvDriveObjectBase__svh
`define GpvDriveObjectBase__svh

virtual class GpvDriveObjectBase extends uvm_object; // {

	function new(string name="GpvDriveObjectBase");
		super.new(name);
	endfunction

endclass // }

`endif
