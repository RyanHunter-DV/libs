`ifndef rhGpvTypes__svh
`define rhGpvTypes__svh

typedef struct {
	int s;
	int e;
}RhGpvSigPos_t;

`endif
